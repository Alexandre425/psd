package common is
    type alu_operation is (ALU_ADD, ALU_MULT, ALU_OR, ALU_RTR);
end common;