library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package common is
    type complex_matrix is array (7 downto 0) of std_logic_vector(11 downto 0);
end common;
